** Profile: "SCHEMATIC1-Lab1_1.1"  [ D:\KMITL\YEAR1\term2\Circuit&Electronics\Lab1\lab1_1.1-SCHEMATIC1-Lab1_1.1.sim ] 

** Creating circuit file "lab1_1.1-SCHEMATIC1-Lab1_1.1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\Orcad_9.2.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ns 0 1 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\lab1_1.1-SCHEMATIC1.net" 


.END
