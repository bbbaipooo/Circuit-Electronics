** Profile: "SCHEMATIC1-Lab1_1.10"  [ D:\KMITL\year1\term2\Circuit&Electronics\Lab1\lab1_1.9-schematic1-lab1_1.10.sim ] 

** Creating circuit file "lab1_1.9-schematic1-lab1_1.10.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\Orcad_9.2.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 0.1m 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\lab1_1.9-SCHEMATIC1.net" 


.END
