** Profile: "SCHEMATIC1-LAB11-1"  [ D:\KMITL\year1\term2\Circuit&Electronics\LAB\lab11-1-SCHEMATIC1-LAB11-1.sim ] 

** Creating circuit file "lab11-1-SCHEMATIC1-LAB11-1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\Orcad_9.2.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10s 0 0.01m 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\lab11-1-SCHEMATIC1.net" 


.END
