** Profile: "SCHEMATIC1-TEST"  [ D:\KMITL\year1\term2\Circuit&Electronics\test-SCHEMATIC1-TEST.sim ] 

** Creating circuit file "test-SCHEMATIC1-TEST.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\Orcad_9.2.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\test-SCHEMATIC1.net" 


.END
