** Profile: "SCHEMATIC1-Lab1_1.5"  [ D:\KMITL\year1\term2\Circuit&Electronics\Lab1\lab1_1.5-schematic1-lab1_1.5.sim ] 

** Creating circuit file "lab1_1.5-schematic1-lab1_1.5.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\Orcad_9.2.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 10us 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\lab1_1.5-SCHEMATIC1.net" 


.END
