** Profile: "SCHEMATIC1-LAB11-2"  [ D:\KMITL\year1\term2\Circuit&Electronics\LAB\lab11-2-SCHEMATIC1-LAB11-2.sim ] 

** Creating circuit file "lab11-2-SCHEMATIC1-LAB11-2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\Orcad_9.2.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 50ms 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\lab11-2-SCHEMATIC1.net" 


.END
